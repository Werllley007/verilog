module exec01_tb;
    localparam WIDTH
    
endmodule